// top file

module top ()

endmodule
```